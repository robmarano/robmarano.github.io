`ifndef REGISTER_FILE
`define REGISTER_FILE

`include "register.sv"

module register_file
    #(
    parameter DEPTH = 8,  // Number of registers (default 8)
    parameter WIDTH = 8   // Width of each register (inherited or specified)
    ) (
    input logic clk,
    input logic rst,
    input logic enable,

    input logic [$clog2(DEPTH)-1:0] write_addr, // Write address
    input logic [WIDTH-1:0] write_data,      // Write data
    input logic write_en,                  // Write enable
    input logic [$clog2(DEPTH)-1:0] read_addr, // Read address
    output logic [WIDTH-1:0] read_data     // Read data
);

    // Array of registers
    register #( .WIDTH(WIDTH) ) registers [DEPTH-1:0]; // Parameterized register instances

    parameter bit [WIDTH-1:0] ZERO  = '0;

    genvar i;
    generate
        for (i = 0; i < DEPTH; i++) begin
            register #( .WIDTH(WIDTH) ) registers (
                .clk(clk),
                .rst(rst),
                .enable(enable && write_en && (write_addr == i)), // Simplified enable logic
                .d(write_data),
                .q() // Output not directly connected within the array
            );  
        end
    endgenerate
                // .enable(enable),
                // .d( (write_en && (write_addr == i)) ? write_data : ZERO ), // Conditional write

    logic [WIDTH-1:0] read_data_internal; // Intermediate signal
    always_ff @(posedge clk) begin
        read_data_internal <= registers[read_addr].q; // Indexing with read_addr
    end
endmodule

`endif